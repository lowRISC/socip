// See LICENSE for license details.

module nasti_channel_slicer
  #(
    N_PORT = 1                 // number of nasti ports to be sliced, maximal 8
    )
   (
    nasti_channel.slave master,
    nasti_channel.master slave_0, slave_1, slave_2, slave_3, slave_4, slave_5, slave_6, slave_7
    );

   // much easier if Vivado support array of interfaces
   generate
      if(N_PORT > 0) begin
         assign slave_0.aw_id      = master.aw_id[0];
         assign slave_0.aw_addr    = master.aw_addr[0];
         assign slave_0.aw_len     = master.aw_len[0];
         assign slave_0.aw_size    = master.aw_size[0];
         assign slave_0.aw_burst   = master.aw_burst[0];
         assign slave_0.aw_lock    = master.aw_lock[0];
         assign slave_0.aw_cache   = master.aw_cache[0];
         assign slave_0.aw_prot    = master.aw_prot[0];
         assign slave_0.aw_qos     = master.aw_qos[0];
         assign slave_0.aw_region  = master.aw_region[0];
         assign slave_0.aw_user    = master.aw_user[0];
         assign slave_0.aw_valid   = master.aw_valid[0];
         assign slave_0.ar_id      = master.ar_id[0];
         assign slave_0.ar_addr    = master.ar_addr[0];
         assign slave_0.ar_len     = master.ar_len[0];
         assign slave_0.ar_size    = master.ar_size[0];
         assign slave_0.ar_burst   = master.ar_burst[0];
         assign slave_0.ar_lock    = master.ar_lock[0];
         assign slave_0.ar_cache   = master.ar_cache[0];
         assign slave_0.ar_prot    = master.ar_prot[0];
         assign slave_0.ar_qos     = master.ar_qos[0];
         assign slave_0.ar_region  = master.ar_region[0];
         assign slave_0.ar_user    = master.ar_user[0];
         assign slave_0.ar_valid   = master.ar_valid[0];
         assign slave_0.w_data     = master.w_data[0];
         assign slave_0.w_strb     = master.w_strb[0];
         assign slave_0.w_last     = master.w_last[0];
         assign slave_0.w_user     = master.w_user[0];
         assign slave_0.w_valid    = master.w_valid[0];
         assign slave_0.b_ready    = master.b_ready[0];
         assign slave_0.r_ready    = master.r_ready[0];
         assign master.aw_ready[0] = slave_0.aw_ready;
         assign master.ar_ready[0] = slave_0.ar_ready;
         assign master.w_ready[0]  = slave_0.w_ready;
         assign master.b_id[0]     = slave_0.b_id;
         assign master.b_resp[0]   = slave_0.b_resp;
         assign master.b_user[0]   = slave_0.b_user;
         assign master.b_valid[0]  = slave_0.b_valid;
         assign master.r_data[0]   = slave_0.r_data;
         assign master.r_last[0]   = slave_0.r_last;
         assign master.r_id[0]     = slave_0.r_id;
         assign master.r_resp[0]   = slave_0.r_resp;
         assign master.r_user[0]   = slave_0.r_user;
         assign master.r_valid[0]  = slave_0.r_valid;
      end

      if(N_PORT > 1) begin
         assign slave_1.aw_id      = master.aw_id[1];
         assign slave_1.aw_addr    = master.aw_addr[1];
         assign slave_1.aw_len     = master.aw_len[1];
         assign slave_1.aw_size    = master.aw_size[1];
         assign slave_1.aw_burst   = master.aw_burst[1];
         assign slave_1.aw_lock    = master.aw_lock[1];
         assign slave_1.aw_cache   = master.aw_cache[1];
         assign slave_1.aw_prot    = master.aw_prot[1];
         assign slave_1.aw_qos     = master.aw_qos[1];
         assign slave_1.aw_region  = master.aw_region[1];
         assign slave_1.aw_user    = master.aw_user[1];
         assign slave_1.aw_valid   = master.aw_valid[1];
         assign slave_1.ar_id      = master.ar_id[1];
         assign slave_1.ar_addr    = master.ar_addr[1];
         assign slave_1.ar_len     = master.ar_len[1];
         assign slave_1.ar_size    = master.ar_size[1];
         assign slave_1.ar_burst   = master.ar_burst[1];
         assign slave_1.ar_lock    = master.ar_lock[1];
         assign slave_1.ar_cache   = master.ar_cache[1];
         assign slave_1.ar_prot    = master.ar_prot[1];
         assign slave_1.ar_qos     = master.ar_qos[1];
         assign slave_1.ar_region  = master.ar_region[1];
         assign slave_1.ar_user    = master.ar_user[1];
         assign slave_1.ar_valid   = master.ar_valid[1];
         assign slave_1.w_data     = master.w_data[1];
         assign slave_1.w_strb     = master.w_strb[1];
         assign slave_1.w_last     = master.w_last[1];
         assign slave_1.w_user     = master.w_user[1];
         assign slave_1.w_valid    = master.w_valid[1];
         assign slave_1.b_ready    = master.b_ready[1];
         assign slave_1.r_ready    = master.r_ready[1];
         assign master.aw_ready[1] = slave_1.aw_ready;
         assign master.ar_ready[1] = slave_1.ar_ready;
         assign master.w_ready[1]  = slave_1.w_ready;
         assign master.b_id[1]     = slave_1.b_id;
         assign master.b_resp[1]   = slave_1.b_resp;
         assign master.b_user[1]   = slave_1.b_user;
         assign master.b_valid[1]  = slave_1.b_valid;
         assign master.r_data[1]   = slave_1.r_data;
         assign master.r_last[1]   = slave_1.r_last;
         assign master.r_id[1]     = slave_1.r_id;
         assign master.r_resp[1]   = slave_1.r_resp;
         assign master.r_user[1]   = slave_1.r_user;
         assign master.r_valid[1]  = slave_1.r_valid;
      end

      if(N_PORT > 2) begin
         assign slave_2.aw_id      = master.aw_id[2];
         assign slave_2.aw_addr    = master.aw_addr[2];
         assign slave_2.aw_len     = master.aw_len[2];
         assign slave_2.aw_size    = master.aw_size[2];
         assign slave_2.aw_burst   = master.aw_burst[2];
         assign slave_2.aw_lock    = master.aw_lock[2];
         assign slave_2.aw_cache   = master.aw_cache[2];
         assign slave_2.aw_prot    = master.aw_prot[2];
         assign slave_2.aw_qos     = master.aw_qos[2];
         assign slave_2.aw_region  = master.aw_region[2];
         assign slave_2.aw_user    = master.aw_user[2];
         assign slave_2.aw_valid   = master.aw_valid[2];
         assign slave_2.ar_id      = master.ar_id[2];
         assign slave_2.ar_addr    = master.ar_addr[2];
         assign slave_2.ar_len     = master.ar_len[2];
         assign slave_2.ar_size    = master.ar_size[2];
         assign slave_2.ar_burst   = master.ar_burst[2];
         assign slave_2.ar_lock    = master.ar_lock[2];
         assign slave_2.ar_cache   = master.ar_cache[2];
         assign slave_2.ar_prot    = master.ar_prot[2];
         assign slave_2.ar_qos     = master.ar_qos[2];
         assign slave_2.ar_region  = master.ar_region[2];
         assign slave_2.ar_user    = master.ar_user[2];
         assign slave_2.ar_valid   = master.ar_valid[2];
         assign slave_2.w_data     = master.w_data[2];
         assign slave_2.w_strb     = master.w_strb[2];
         assign slave_2.w_last     = master.w_last[2];
         assign slave_2.w_user     = master.w_user[2];
         assign slave_2.w_valid    = master.w_valid[2];
         assign slave_2.b_ready    = master.b_ready[2];
         assign slave_2.r_ready    = master.r_ready[2];
         assign master.aw_ready[2] = slave_2.aw_ready;
         assign master.ar_ready[2] = slave_2.ar_ready;
         assign master.w_ready[2]  = slave_2.w_ready;
         assign master.b_id[2]     = slave_2.b_id;
         assign master.b_resp[2]   = slave_2.b_resp;
         assign master.b_user[2]   = slave_2.b_user;
         assign master.b_valid[2]  = slave_2.b_valid;
         assign master.r_data[2]   = slave_2.r_data;
         assign master.r_last[2]   = slave_2.r_last;
         assign master.r_id[2]     = slave_2.r_id;
         assign master.r_resp[2]   = slave_2.r_resp;
         assign master.r_user[2]   = slave_2.r_user;
         assign master.r_valid[2]  = slave_2.r_valid;
      end

      if(N_PORT > 3) begin
         assign slave_3.aw_id      = master.aw_id[3];
         assign slave_3.aw_addr    = master.aw_addr[3];
         assign slave_3.aw_len     = master.aw_len[3];
         assign slave_3.aw_size    = master.aw_size[3];
         assign slave_3.aw_burst   = master.aw_burst[3];
         assign slave_3.aw_lock    = master.aw_lock[3];
         assign slave_3.aw_cache   = master.aw_cache[3];
         assign slave_3.aw_prot    = master.aw_prot[3];
         assign slave_3.aw_qos     = master.aw_qos[3];
         assign slave_3.aw_region  = master.aw_region[3];
         assign slave_3.aw_user    = master.aw_user[3];
         assign slave_3.aw_valid   = master.aw_valid[3];
         assign slave_3.ar_id      = master.ar_id[3];
         assign slave_3.ar_addr    = master.ar_addr[3];
         assign slave_3.ar_len     = master.ar_len[3];
         assign slave_3.ar_size    = master.ar_size[3];
         assign slave_3.ar_burst   = master.ar_burst[3];
         assign slave_3.ar_lock    = master.ar_lock[3];
         assign slave_3.ar_cache   = master.ar_cache[3];
         assign slave_3.ar_prot    = master.ar_prot[3];
         assign slave_3.ar_qos     = master.ar_qos[3];
         assign slave_3.ar_region  = master.ar_region[3];
         assign slave_3.ar_user    = master.ar_user[3];
         assign slave_3.ar_valid   = master.ar_valid[3];
         assign slave_3.w_data     = master.w_data[3];
         assign slave_3.w_strb     = master.w_strb[3];
         assign slave_3.w_last     = master.w_last[3];
         assign slave_3.w_user     = master.w_user[3];
         assign slave_3.w_valid    = master.w_valid[3];
         assign slave_3.b_ready    = master.b_ready[3];
         assign slave_3.r_ready    = master.r_ready[3];
         assign master.aw_ready[3] = slave_3.aw_ready;
         assign master.ar_ready[3] = slave_3.ar_ready;
         assign master.w_ready[3]  = slave_3.w_ready;
         assign master.b_id[3]     = slave_3.b_id;
         assign master.b_resp[3]   = slave_3.b_resp;
         assign master.b_user[3]   = slave_3.b_user;
         assign master.b_valid[3]  = slave_3.b_valid;
         assign master.r_data[3]   = slave_3.r_data;
         assign master.r_last[3]   = slave_3.r_last;
         assign master.r_id[3]     = slave_3.r_id;
         assign master.r_resp[3]   = slave_3.r_resp;
         assign master.r_user[3]   = slave_3.r_user;
         assign master.r_valid[3]  = slave_3.r_valid;
      end

      if(N_PORT > 4) begin
         assign slave_4.aw_id      = master.aw_id[4];
         assign slave_4.aw_addr    = master.aw_addr[4];
         assign slave_4.aw_len     = master.aw_len[4];
         assign slave_4.aw_size    = master.aw_size[4];
         assign slave_4.aw_burst   = master.aw_burst[4];
         assign slave_4.aw_lock    = master.aw_lock[4];
         assign slave_4.aw_cache   = master.aw_cache[4];
         assign slave_4.aw_prot    = master.aw_prot[4];
         assign slave_4.aw_qos     = master.aw_qos[4];
         assign slave_4.aw_region  = master.aw_region[4];
         assign slave_4.aw_user    = master.aw_user[4];
         assign slave_4.aw_valid   = master.aw_valid[4];
         assign slave_4.ar_id      = master.ar_id[4];
         assign slave_4.ar_addr    = master.ar_addr[4];
         assign slave_4.ar_len     = master.ar_len[4];
         assign slave_4.ar_size    = master.ar_size[4];
         assign slave_4.ar_burst   = master.ar_burst[4];
         assign slave_4.ar_lock    = master.ar_lock[4];
         assign slave_4.ar_cache   = master.ar_cache[4];
         assign slave_4.ar_prot    = master.ar_prot[4];
         assign slave_4.ar_qos     = master.ar_qos[4];
         assign slave_4.ar_region  = master.ar_region[4];
         assign slave_4.ar_user    = master.ar_user[4];
         assign slave_4.ar_valid   = master.ar_valid[4];
         assign slave_4.w_data     = master.w_data[4];
         assign slave_4.w_strb     = master.w_strb[4];
         assign slave_4.w_last     = master.w_last[4];
         assign slave_4.w_user     = master.w_user[4];
         assign slave_4.w_valid    = master.w_valid[4];
         assign slave_4.b_ready    = master.b_ready[4];
         assign slave_4.r_ready    = master.r_ready[4];
         assign master.aw_ready[4] = slave_4.aw_ready;
         assign master.ar_ready[4] = slave_4.ar_ready;
         assign master.w_ready[4]  = slave_4.w_ready;
         assign master.b_id[4]     = slave_4.b_id;
         assign master.b_resp[4]   = slave_4.b_resp;
         assign master.b_user[4]   = slave_4.b_user;
         assign master.b_valid[4]  = slave_4.b_valid;
         assign master.r_data[4]   = slave_4.r_data;
         assign master.r_last[4]   = slave_4.r_last;
         assign master.r_id[4]     = slave_4.r_id;
         assign master.r_resp[4]   = slave_4.r_resp;
         assign master.r_user[4]   = slave_4.r_user;
         assign master.r_valid[4]  = slave_4.r_valid;
      end

      if(N_PORT > 5) begin
         assign slave_5.aw_id      = master.aw_id[5];
         assign slave_5.aw_addr    = master.aw_addr[5];
         assign slave_5.aw_len     = master.aw_len[5];
         assign slave_5.aw_size    = master.aw_size[5];
         assign slave_5.aw_burst   = master.aw_burst[5];
         assign slave_5.aw_lock    = master.aw_lock[5];
         assign slave_5.aw_cache   = master.aw_cache[5];
         assign slave_5.aw_prot    = master.aw_prot[5];
         assign slave_5.aw_qos     = master.aw_qos[5];
         assign slave_5.aw_region  = master.aw_region[5];
         assign slave_5.aw_user    = master.aw_user[5];
         assign slave_5.aw_valid   = master.aw_valid[5];
         assign slave_5.ar_id      = master.ar_id[5];
         assign slave_5.ar_addr    = master.ar_addr[5];
         assign slave_5.ar_len     = master.ar_len[5];
         assign slave_5.ar_size    = master.ar_size[5];
         assign slave_5.ar_burst   = master.ar_burst[5];
         assign slave_5.ar_lock    = master.ar_lock[5];
         assign slave_5.ar_cache   = master.ar_cache[5];
         assign slave_5.ar_prot    = master.ar_prot[5];
         assign slave_5.ar_qos     = master.ar_qos[5];
         assign slave_5.ar_region  = master.ar_region[5];
         assign slave_5.ar_user    = master.ar_user[5];
         assign slave_5.ar_valid   = master.ar_valid[5];
         assign slave_5.w_data     = master.w_data[5];
         assign slave_5.w_strb     = master.w_strb[5];
         assign slave_5.w_last     = master.w_last[5];
         assign slave_5.w_user     = master.w_user[5];
         assign slave_5.w_valid    = master.w_valid[5];
         assign slave_5.b_ready    = master.b_ready[5];
         assign slave_5.r_ready    = master.r_ready[5];
         assign master.aw_ready[5] = slave_5.aw_ready;
         assign master.ar_ready[5] = slave_5.ar_ready;
         assign master.w_ready[5]  = slave_5.w_ready;
         assign master.b_id[5]     = slave_5.b_id;
         assign master.b_resp[5]   = slave_5.b_resp;
         assign master.b_user[5]   = slave_5.b_user;
         assign master.b_valid[5]  = slave_5.b_valid;
         assign master.r_data[5]   = slave_5.r_data;
         assign master.r_last[5]   = slave_5.r_last;
         assign master.r_id[5]     = slave_5.r_id;
         assign master.r_resp[5]   = slave_5.r_resp;
         assign master.r_user[5]   = slave_5.r_user;
         assign master.r_valid[5]  = slave_5.r_valid;
      end

      if(N_PORT > 6) begin
         assign slave_6.aw_id      = master.aw_id[6];
         assign slave_6.aw_addr    = master.aw_addr[6];
         assign slave_6.aw_len     = master.aw_len[6];
         assign slave_6.aw_size    = master.aw_size[6];
         assign slave_6.aw_burst   = master.aw_burst[6];
         assign slave_6.aw_lock    = master.aw_lock[6];
         assign slave_6.aw_cache   = master.aw_cache[6];
         assign slave_6.aw_prot    = master.aw_prot[6];
         assign slave_6.aw_qos     = master.aw_qos[6];
         assign slave_6.aw_region  = master.aw_region[6];
         assign slave_6.aw_user    = master.aw_user[6];
         assign slave_6.aw_valid   = master.aw_valid[6];
         assign slave_6.ar_id      = master.ar_id[6];
         assign slave_6.ar_addr    = master.ar_addr[6];
         assign slave_6.ar_len     = master.ar_len[6];
         assign slave_6.ar_size    = master.ar_size[6];
         assign slave_6.ar_burst   = master.ar_burst[6];
         assign slave_6.ar_lock    = master.ar_lock[6];
         assign slave_6.ar_cache   = master.ar_cache[6];
         assign slave_6.ar_prot    = master.ar_prot[6];
         assign slave_6.ar_qos     = master.ar_qos[6];
         assign slave_6.ar_region  = master.ar_region[6];
         assign slave_6.ar_user    = master.ar_user[6];
         assign slave_6.ar_valid   = master.ar_valid[6];
         assign slave_6.w_data     = master.w_data[6];
         assign slave_6.w_strb     = master.w_strb[6];
         assign slave_6.w_last     = master.w_last[6];
         assign slave_6.w_user     = master.w_user[6];
         assign slave_6.w_valid    = master.w_valid[6];
         assign slave_6.b_ready    = master.b_ready[6];
         assign slave_6.r_ready    = master.r_ready[6];
         assign master.aw_ready[6] = slave_6.aw_ready;
         assign master.ar_ready[6] = slave_6.ar_ready;
         assign master.w_ready[6]  = slave_6.w_ready;
         assign master.b_id[6]     = slave_6.b_id;
         assign master.b_resp[6]   = slave_6.b_resp;
         assign master.b_user[6]   = slave_6.b_user;
         assign master.b_valid[6]  = slave_6.b_valid;
         assign master.r_data[6]   = slave_6.r_data;
         assign master.r_last[6]   = slave_6.r_last;
         assign master.r_id[6]     = slave_6.r_id;
         assign master.r_resp[6]   = slave_6.r_resp;
         assign master.r_user[6]   = slave_6.r_user;
         assign master.r_valid[6]  = slave_6.r_valid;
      end

      if(N_PORT > 7) begin
         assign slave_7.aw_id      = master.aw_id[7];
         assign slave_7.aw_addr    = master.aw_addr[7];
         assign slave_7.aw_len     = master.aw_len[7];
         assign slave_7.aw_size    = master.aw_size[7];
         assign slave_7.aw_burst   = master.aw_burst[7];
         assign slave_7.aw_lock    = master.aw_lock[7];
         assign slave_7.aw_cache   = master.aw_cache[7];
         assign slave_7.aw_prot    = master.aw_prot[7];
         assign slave_7.aw_qos     = master.aw_qos[7];
         assign slave_7.aw_region  = master.aw_region[7];
         assign slave_7.aw_user    = master.aw_user[7];
         assign slave_7.aw_valid   = master.aw_valid[7];
         assign slave_7.ar_id      = master.ar_id[7];
         assign slave_7.ar_addr    = master.ar_addr[7];
         assign slave_7.ar_len     = master.ar_len[7];
         assign slave_7.ar_size    = master.ar_size[7];
         assign slave_7.ar_burst   = master.ar_burst[7];
         assign slave_7.ar_lock    = master.ar_lock[7];
         assign slave_7.ar_cache   = master.ar_cache[7];
         assign slave_7.ar_prot    = master.ar_prot[7];
         assign slave_7.ar_qos     = master.ar_qos[7];
         assign slave_7.ar_region  = master.ar_region[7];
         assign slave_7.ar_user    = master.ar_user[7];
         assign slave_7.ar_valid   = master.ar_valid[7];
         assign slave_7.w_data     = master.w_data[7];
         assign slave_7.w_strb     = master.w_strb[7];
         assign slave_7.w_last     = master.w_last[7];
         assign slave_7.w_user     = master.w_user[7];
         assign slave_7.w_valid    = master.w_valid[7];
         assign slave_7.b_ready    = master.b_ready[7];
         assign slave_7.r_ready    = master.r_ready[7];
         assign master.aw_ready[7] = slave_7.aw_ready;
         assign master.ar_ready[7] = slave_7.ar_ready;
         assign master.w_ready[7]  = slave_7.w_ready;
         assign master.b_id[7]     = slave_7.b_id;
         assign master.b_resp[7]   = slave_7.b_resp;
         assign master.b_user[7]   = slave_7.b_user;
         assign master.b_valid[7]  = slave_7.b_valid;
         assign master.r_data[7]   = slave_7.r_data;
         assign master.r_last[7]   = slave_7.r_last;
         assign master.r_id[7]     = slave_7.r_id;
         assign master.r_resp[7]   = slave_7.r_resp;
         assign master.r_user[7]   = slave_7.r_user;
         assign master.r_valid[7]  = slave_7.r_valid;
      end
   endgenerate

endmodule // nasti_channel_slicer
